-- }}}                                                                                                    
begin                                                                                                         

   --! @brief DUT Port Map                                                                                   
   -- {{{                  
