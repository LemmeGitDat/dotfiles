library ieee;                                                                                                 
use ieee.std_logic_1164.all;                                                                                  

--! Entity Declaration                                                                                        
-- {{{                                                                                                        
entity tb_template is                                                                                         
   end tb_template;                                                                                           
-- }}}                                                                                                        

--! @brief Architecture Description                                                                           
-- {{{                                                                                                        
architecture arch of tb_template is                                                                           
   --! @brief Signal Declarations                                                                            
   -- {{{                                                                                                    
   constant clk_period : time := 100 ns;    
